module hex_digits(
  input       clk_i, rst_i
  input [4:0] hex0,     // Входной сигнал со значением цифры, выводимой на нулевой (самый правый) индикатор
  input [4:0] hex1,     // Входной сигнал со значением цифры, выводимой на первый индикатор
  input [4:0] hex2,     // Входной сигнал со значением цифры, выводимой на второй индикатор
  input [4:0] hex3,     // Входной сигнал со значением цифры, выводимой на третий индикатор
  input [4:0] hex4,     // Входной сигнал со значением цифры, выводимой на четвертый индикатор
  input [4:0] hex5,     // Входной сигнал со значением цифры, выводимой на пятый индикатор
  input [4:0] hex6,     // Входной сигнал со значением цифры, выводимой на шестой индикатор
  input [4:0] hex7,     // Входной сигнал со значением цифры, выводимой на седьмой индикатор

  output [6:0] hex_led  // Выходной сигнал, контролирующий каждый отдельный светодиод индикатора
  output [7:0] hex_sel  // Выходной сигнал, указывающий на какой индикатор выставляется hex_led
);
endmodule